library verilog;
use verilog.vl_types.all;
entity lab2part2_vlg_vec_tst is
end lab2part2_vlg_vec_tst;

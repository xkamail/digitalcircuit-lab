library verilog;
use verilog.vl_types.all;
entity lab2part6_vlg_vec_tst is
end lab2part6_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity lab3part3_vlg_vec_tst is
end lab3part3_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity lab4part5_vlg_vec_tst is
end lab4part5_vlg_vec_tst;

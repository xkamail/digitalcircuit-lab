library verilog;
use verilog.vl_types.all;
entity lab7part4_vlg_vec_tst is
end lab7part4_vlg_vec_tst;

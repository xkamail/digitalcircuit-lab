library verilog;
use verilog.vl_types.all;
entity lab5part3_vlg_vec_tst is
end lab5part3_vlg_vec_tst;

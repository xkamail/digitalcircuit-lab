library verilog;
use verilog.vl_types.all;
entity lab3part4_vlg_vec_tst is
end lab3part4_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity lab1part4_vlg_sample_tst is
    port(
        c0              : in     vl_logic;
        c1              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end lab1part4_vlg_sample_tst;

library verilog;
use verilog.vl_types.all;
entity lab4part1_vlg_vec_tst is
end lab4part1_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity lab4part3_vlg_sample_tst is
    port(
        clock50         : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end lab4part3_vlg_sample_tst;

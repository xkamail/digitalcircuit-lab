library verilog;
use verilog.vl_types.all;
entity lab4part4_vlg_vec_tst is
end lab4part4_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity lab2part5_vlg_vec_tst is
end lab2part5_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity lab8part1_vlg_vec_tst is
end lab8part1_vlg_vec_tst;

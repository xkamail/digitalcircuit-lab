library verilog;
use verilog.vl_types.all;
entity lab5part1_vlg_vec_tst is
end lab5part1_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity lab5part1_vlg_sample_tst is
    port(
        key0            : in     vl_logic;
        reset           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end lab5part1_vlg_sample_tst;

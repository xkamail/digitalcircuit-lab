library verilog;
use verilog.vl_types.all;
entity lab3part3 is
    port(
        D               : in     vl_logic;
        Clk             : in     vl_logic;
        Q               : out    vl_logic
    );
end lab3part3;

library verilog;
use verilog.vl_types.all;
entity lab1part2_vlg_vec_tst is
end lab1part2_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity lab5part2_vlg_vec_tst is
end lab5part2_vlg_vec_tst;

library ieee;
use ieee.std_logic_1164.all;

entity every_seconds is
	port (
		clock50 : in std_logic;
		
	);
end every_seconds;
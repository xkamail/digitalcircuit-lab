library verilog;
use verilog.vl_types.all;
entity lab6part4_vlg_vec_tst is
end lab6part4_vlg_vec_tst;

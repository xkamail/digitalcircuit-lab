library verilog;
use verilog.vl_types.all;
entity lab3part5_vlg_vec_tst is
end lab3part5_vlg_vec_tst;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity decimal_encoder is 
	port (
		x : std_logic_vector(6 downto 0)
	);
end decimal_encoder;
architecture bhv of decimal_encoder is

begin

end bhv;
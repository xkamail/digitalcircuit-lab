library verilog;
use verilog.vl_types.all;
entity lab1part3_vlg_check_tst is
    port(
        m               : in     vl_logic_vector(1 downto 0);
        sampler_rx      : in     vl_logic
    );
end lab1part3_vlg_check_tst;

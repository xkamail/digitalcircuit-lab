library verilog;
use verilog.vl_types.all;
entity lab7part3_vlg_vec_tst is
end lab7part3_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity lab3part1_vlg_vec_tst is
end lab3part1_vlg_vec_tst;

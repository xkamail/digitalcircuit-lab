library verilog;
use verilog.vl_types.all;
entity lab3part1 is
    port(
        Clk             : in     vl_logic;
        R               : in     vl_logic;
        S               : in     vl_logic;
        Q               : out    vl_logic
    );
end lab3part1;

library verilog;
use verilog.vl_types.all;
entity lab3part3_vlg_check_tst is
    port(
        Q               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab3part3_vlg_check_tst;
